-- 
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;


ENTITY IR IS
	PORT(
		DATA : IN STD_LOGIC_VECTOR(11 DOWNTO 0);
		CLK : IN STD_LOGIC;
		WREN : IN STD_LOGIC;
		Q : OUT STD_LOGIC_VECTOR(11 DOWNTO 0)
	);
END IR;

ARCHITECTURE SYN OF IR IS
	SIGNAL d : STD_LOGIC_VECTOR(11 DOWNTO 0);
BEGIN
	PROCESS(CLK, WREN)
	BEGIN
		IF CLK'EVENT AND CLK = '1' THEN
			IF WREN = '1' THEN
				d <= DATA;
			END IF;
		END IF;
	END PROCESS;

	Q <= d;

END SYN;
