
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY reg_B IS
	PORT(
		DATA : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		GATE : IN STD_LOGIC;
		Q : OUT STD_LOGIC_VECTOR(5 DOWNTO 0)
	);
END reg_B;

ARCHITECTURE SYN OF reg_B IS
BEGIN
	PROCESS(GATE)
	BEGIN
		IF GATE = '1' THEN
			Q <= DATA;
		END IF;
	END PROCESS;

END SYN;

