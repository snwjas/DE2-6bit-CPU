-- 

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY comparator IS
	PORT(
		A : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		B : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		Q : OUT STD_LOGIC
	);
END comparator;

ARCHITECTURE SYN OF comparator IS
BEGIN
	Q <= '1' WHEN A = B ELSE '0';
END SYN;