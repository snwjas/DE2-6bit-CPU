
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY PM IS
	PORT (
		DATA: IN STD_LOGIC_VECTOR(11 DOWNTO 0);
		WCLK: IN STD_LOGIC;
		WADR: IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		RCLK: IN STD_LOGIC;
		RADR: IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		Q: OUT STD_LOGIC_VECTOR(11 DOWNTO 0)
	);
END PM;

ARCHITECTURE SYN OF PM IS
	-- row
	TYPE MEM IS ARRAY(0 TO 15) OF
	-- col
	STD_LOGIC_VECTOR(11 DOWNTO 0);
	SIGNAL RAMTMP: MEM;
BEGIN
	WR: PROCESS(WCLK)
	BEGIN
		IF WCLK'EVENT AND WCLK = '1' THEN
			RAMTMP(CONV_INTEGER(WADR)) <= DATA;
		END IF;
	END PROCESS;

	RD: PROCESS(RCLK)
	BEGIN
		IF RCLK'EVENT AND RCLK = '1' THEN
			Q <= RAMTMP(CONV_INTEGER(RADR));
		END IF;
	END PROCESS;
END SYN;